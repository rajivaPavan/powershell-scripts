library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity template is
    -- port();
end template;

architecture Behavioral of template is

begin

end Behavioral;
